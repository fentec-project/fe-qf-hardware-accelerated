`timescale	1ns/1ps
///////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////
module maab
	(
	clk,
	a,
	b,
	c,
	d,
	p
	);

	// Ports ///////////////////////////////////////////////////////////////////
	input			clk;

	input	[63:0]	a;
	input	[63:0]	b;
	input	[63:0]	c;
	input	[63:0]	d;

	output	[127:0]	p;

	// Internal signal and register ////////////////////////////////////////////
	wire	[64:0] 	w11;
	wire	[63:0] 	w12;
	wire	[32:0] 	w13;
	wire	[32:0] 	w14;
	wire	[63:0] 	w15;

	reg		[64:0]	r11;
	reg		[63:0]	r12;
	reg		[32:0]	r13;
	reg		[32:0]	r14;
	reg		[63:0]	r15;

	wire	[65:0] 	w21;
	wire	[65:0] 	w22;
	wire	[64:0] 	w23;

	reg		[65:0]	r21;
	reg		[65:0]	r22;
	reg		[64:0]	r23;
	reg		[63:0]	r24;

	wire	[32:0] 	w31;
	wire	[65:0] 	w32;
	wire	[95:0] 	w33;

	reg		[31:0]	r31;
	reg		[1:0]	r32;
	reg		[31:0]	r33;
	reg				r34;
	reg		[63:0]	r35;
	reg		[63:0]	r36;

	// Assignments //////////////////////////////////////////////////////////////
	assign w11 = c + d;
	assign w12 = a[31:0] * b[31:0];
	assign w13 = b[63:32] + b[31:0];
	assign w14 = a[63:32] + a[31:0];
	assign w15 = a[63:32] * b[63:32];

	assign w21 = r11 + r12;
	assign w22 = r13 * r14;
	assign w23 = ~(r12 + r15);

	assign w32 = r22 + {1'b1, r23} + 1'b1;
	assign w33 = {w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65],
				  w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], 
				  w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], 
				  w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:0]};
	assign w31 = w33[31:0] + r21[63:32];

	assign p[31:0] = r31;
	assign p[63:32] = r33;
	assign p[127:64] = r32 + r34 + r35 + r36;

	// Sequential procedures ///////////////////////////////////////////////////
	always @(posedge clk)
	begin
		r11 <= w11;
		r12 <= w12;
		r13 <= w13;
		r14 <= w14;
		r15 <= w15;
	end
	
	always @(posedge clk)
	begin
		r21 <= w21;
		r22 <= w22;
		r23 <= w23;
		r24 <= r15;
	end
	
	always @(posedge clk)
	begin
		r31 <= r21[31:0];
		r32 <= r21[65:64];
		r33 <= w31[31:0];
		r34 <= w31[32:32];
		r35 <= w33[95:32];
		r36 <= r24;
	end

	////////////////////////////////////////////////////////////////////////////
endmodule

/*///////////////////////////////////////////////////////////////////////////////
module maab
	(
	clk,
	a,
	b,
	c,
	d,
	p
	);

	// Ports ///////////////////////////////////////////////////////////////////
	input			clk;

	input	[63:0]	a;
	input	[63:0]	b;
	input	[63:0]	c;
	input	[63:0]	d;

	output	[127:0]	p;

	// Internal signal and register ////////////////////////////////////////////
	wire	[64:0] 	w11;
	wire	[63:0] 	w12;
	wire	[32:0] 	w13;
	wire	[32:0] 	w14;
	wire	[63:0] 	w15;

	reg		[64:0]	r11;
	reg		[32:0]	r13;
	reg		[32:0]	r14;

	wire	[65:0] 	w21;
	wire	[65:0] 	w22;
	wire	[64:0] 	w23;

	reg		[65:0]	r21;
	reg		[64:0]	r23;
	reg		[63:0]	r24;

	wire	[32:0] 	w31;
	wire	[65:0] 	w32;
	wire	[95:0] 	w33;

	reg		[31:0]	r31;
	reg		[1:0]	r32;
	reg		[31:0]	r33;
	reg				r34;
	reg		[63:0]	r35;
	reg		[63:0]	r36;

	// Assignments //////////////////////////////////////////////////////////////
	assign w11 = c + d;
	assign w13 = b[63:32] + b[31:0];
	assign w14 = a[63:32] + a[31:0];

	assign w21 = r11 + w12;
	assign w23 = ~(w12 + w15);

	assign w32 = w22 + {1'b1, r23} + 1'b1;
	assign w33 = {w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65],
				  w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], 
				  w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], 
				  w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:65], w32[65:0]};
	assign w31 = w33[31:0] + r21[63:32];

	assign p[31:0] = r31;
	assign p[63:32] = r33;
	assign p[127:64] = r32 + r34 + r35 + r36;

	// Sequential procedures ///////////////////////////////////////////////////
	always @(posedge clk)
	begin
		r11 <= w11;
		r13 <= w13;
		r14 <= w14;
	end
	
	always @(posedge clk)
	begin
		r21 <= w21;
		r23 <= w23;
		r24 <= w15;
	end
	
	always @(posedge clk)
	begin
		r31 <= r21[31:0];
		r32 <= r21[65:64];
		r33 <= w31[31:0];
		r34 <= w31[32:32];
		r35 <= w33[95:32];
		r36 <= r24;
	end

	////////////////////////////////////////////////////////////////////////////
	mult_32_32_64 mult_32_32_64_u1
	(
	  .clk(clk),
	  .a(a[31:0]),
	  .b(b[31:0]),
	  .p(w12)
	);

	////////////////////////////////////////////////////////////////////////////
	mult_32_32_64 mult_32_32_64_u2
	(
	  .clk(clk),
	  .a(a[63:32]),
	  .b(b[63:32]),
	  .p(w15)
	);

	////////////////////////////////////////////////////////////////////////////
	mult_33_33_66 mult_33_33_66_u1
	(
	  .clk(clk),
	  .a(r13),
	  .b(r14),
	  .p(w22)
	);

	////////////////////////////////////////////////////////////////////////////
endmodule*/
